** Profile: "SCHEMATIC1-OCP"  [ d:\1faculta\onedrive - universitatea politehnica bucuresti\cursuri inregistrate\an 3 sem 1\proiect 1\cad\over current protection\ocp-pspicefiles\schematic1\ocp.sim ] 

** Creating circuit file "OCP.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "D:/OrCAD/OrCAD_16.6_Lite/tools/pspice/library/MJD31CG.lib" 
.LIB "D:/OrCAD/OrCAD_16.6_Lite/tools/pspice/library/BC817-25.lib" 
.LIB "D:/OrCAD/OrCAD_16.6_Lite/tools/pspice/library/BC807-25.lib" 
.LIB "D:/OrCAD/OrCAD_16.6_Lite/tools/pspice/library/BZX84C10.lib" 
.LIB "D:/OrCAD/OrCAD_16.6_Lite/tools/pspice/library/BZX84C5V1.lib" 
.LIB "D:/OrCAD/OrCAD_16.6_Lite/tools/pspice/library/BZX84C2V7.lib" 
.LIB "D:/OrCAD/OrCAD_16.6_Lite/tools/pspice/library/MMBFJ309LT1G.lib" 
* From [PSPICE NETLIST] section of C:\Users\Tudor\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 20s 0 0.1s 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
